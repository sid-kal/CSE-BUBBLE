module instruction_memory( address , instruction );

    input [15:0] address;
    output [31:0] instruction;
    reg [31:0] mem [65535:0];
    initial begin
        // mem[0]=32'b001100_00001_00000_00000_00000_000001;
        // mem[1]=32'b001101_00000_00001_01000_00000_000000;
        // // mem[3]=32'b000000_00010_00001_00000_00000_000000;

        // // mem[0]=32'b000000_00010_00001_00000_00000_000000;
        // // mem[1]=32'b010100_00000_00000_00000_00000_000010;
        // // mem[4]=32'b000001_00101_00100_00011_00000_000000;
        // // mem[5]=32'b000010_01000_00111_00110_00000_000000;
        // // mem[6]=32'b000011_01011_01010_01001_00000_000000;


        // mem[0]=32'b00010010101101010000000000000001;
        // mem[1]=32'b00010001110011100000000000000000;
        // mem[2]=32'b00110010100011110000000000000000;
        // mem[3]=32'b00010010100101000000000000000001;
        // mem[4]=32'b00010001001010010000000000000000;
        // mem[5]=32'b00110001010011110000000000000000;
        // mem[6]=32'b00010001111011110000000000000000;
        // mem[7]=32'b00101001101011110000000010000000;
        // mem[8]=32'b00000001101011011010100000000000;
        // mem[9]=32'b00110000110011010000000000000000;
        // mem[10]=32'b00110000111011010000000000000001;
        // mem[11]=32'b01011101000001100011100000000000;
        // mem[12]=32'b00111100000010000000000000000011;
        // mem[13]=32'b00110100000001110110100000000000;
        // mem[14]=32'b00110100000001100110100000000000;
        // mem[15]=32'b00010001111011110000000000000001;
        // mem[16]=32'b00000110011101000111000000000000;
        // mem[17]=32'b00111111111011111001111111110110;
        // mem[18]=32'b00010001110011100000000000000000;
        // mem[19]=32'b00010001111011110000000000000000;
        // mem[20]=32'b00111111111011101010011111110011;
    

        mem[0]=32'b000100_01110_01110_0000000000000001;
        // mem[0]=32'b000100_01110_01110_0000000000000001;
        // mem[1]=32'b000100_01110_01110_0000000000000011;
        // mem[2]=32'b000100_01110_01110_0000000000000001;
        // mem[3]=32'b000100_01110_01110_0000000000000011;
        // mem[4]=32'b000100_01110_01110_0000000000000001;

        // mem[0]=32'b000100_10101_10101_0000000000000001;
        // mem[1]=32'b000100_01110_01110_0000000000000000;
        // mem[2]=32'b001100_10100_01111_0000000000000000;
        // mem[3]=32'b000100_10100_10100_0000000000000001;
        // mem[4]=32'b000100_01001_01001_0000000000000000;
        // mem[5]=32'b001100_01010_01111_0000000000000000;
        // mem[6]=32'b000100_01111_01111_0000000000000000;
        // mem[7]=32'b001010_01101_01111_00000_00010_000000;
        // mem[8]=32'b000000_01101_01101_10101_00000000000;
        // mem[9]=32'b001100_00110_01101_0000000000000000;
        // mem[10]=32'b001100_00111_01101_0000000000000001;
        // mem[11]=32'b010111_01000_00110_00111_00000_000000;
        // mem[12]=32'b001111_00000_01000_00000_00000000011;
        // mem[13]=32'b001101_00000_00111_01101_00000_000000;
        // mem[14]=32'b001101_00000_00110_01101_00000_000000;
        // mem[15]=32'b000100_01111_01111_0000000000000001;
        // mem[16]=32'b000001_10011_10100_01110_00000_000000;
        // mem[17]=32'b001111_11111_01111_10011_11111_110110;
        // mem[18]=32'b000100_01110_01110_0000000000000000;
        // mem[19]=32'b000100_01111_01111_0000000000000000;
        // mem[20]=32'b001111_11111_01110_10100_11111_110011;

    end
    assign instruction=(address<=65535)?mem[address]:0;


/*

00010010101101010000000000000001
00010001110011100000000000000000
00110010100011110000000000000000
00010010100101000000000000000001
00010001001010010000000000000000
00110001010011110000000000000000
00010001111011110000000000000000
00101001101011110000000010000000
00000001101011011010100000000000
00110000110011010000000000000000
00110000111011010000000000000001
01011101000001100011100000000000
00111100000010000000000000000011
00110100000001110110100000000000
00110100000001100110100000000000
00010001111011110000000000000001
00000110011101000111000000000000
00111111111011111001111111110110
00010001110011100000000000000000
00010001111011110000000000000000
00111111111011101010011111110011

*/


endmodule